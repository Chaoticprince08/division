module non_restoring_division_datapath (
    input clk,
    input rst,
    input [15:0] dividend,
    input [15:0] divisor,
);
    
endmodule